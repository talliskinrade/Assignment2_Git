LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.all;
USE work.common_pack.all;

ENTITY cmdProc IS
    PORT (
        clk: IN std_logic;
        reset: IN std_logic;
        rxNow: IN std_logic; -- Equivalent to RX's dataReady signal
        rxData: IN std_logic_vector (7 downto 0);
        txData: OUT std_logic_vector (7 downto 0);
        rxDone: OUT std_logic;
        ovErr: IN std_logic;
        framErr: IN std_logic;
        txNow: OUT std_logic;
        txDone: IN std_logic;
        start: OUT std_logic;
        numWords_bcd: OUT BCD_ARRAY_TYPE(2 downto 0);
        dataReady: IN std_logic;
        byte: IN std_logic_vector(7 downto 0);
        maxIndex: IN BCD_ARRAY_TYPE(2 downto 0);
        dataResults: IN CHAR_ARRAY_TYPE(0 to RESULT_BYTE_NUM-1);
        seqDone: IN std_logic
    );
END cmdProc;

ARCHITECTURE behavioural OF cmdProc IS
-- State Declaration
-- ALL STATE TYPES
	TYPE state_type IS (
	   INIT,
	   RECEIVE_DATA,
	   ECHO_DATA,
	   CHECK_COMMANDS,
	   RESET_COUNT,
	   INCREMENT_COUNT,
	   BYTE_TO_BCD,
	   SEND_TO_DP,
	   BYTE_TO_ASCII,
	   SET_TX,
	   SEND_TX,
	   STORE_RESULTS,
	   BYTE_TO_ASCII_L,
	   RESET_COUNTER_3,
	   SET_TX_L,
	   SEND_TX_L,
	   BYTE_AND_BCD_TO_ASCII,
	   RESET_COUNTER_6,
	   SET_TX_P,
	   SEND_TX_P,
	   DONE
	);
 
-- Signal Declaration
    SIGNAL cur_state, next_state: state_type;
	SIGNAL counter7: integer range 0 to 7;
	SIGNAL counter3: integer range 0 to 3;
	SIGNAL counterA3: integer range 0 to 3;
	SIGNAL receivedDataFlag, sentDataFlag, byteToBCDFlag: std_logic;
	SIGNAL dataBuffer: std_logic_vector (7 downto 0) := "11111111";
	SIGNAL numWordsBuffer: std_logic_vector (11 downto 0) := "000000000000";
	
-------------------------------------------------------------------
--Component Instantiation

--    COMPONENT terminal_echo
--    PORT (
--        clk: IN STD_LOGIC;
--        reset: IN STD_LOGIC;
--        rxNow: IN STD_LOGIC;
--        txDone: IN STD_LOGIC;
--        rxData: IN STD_LOGIC_VECTOR (7 downto 0);
--        txData: OUT STD_LOGIC_VECTOR (7 downto 0);
--        txNow: OUT STD_LOGIC;
--        rxDone: OUT STD_LOGIC
--    );
--    END COMPONENT;
    
--    FOR behavTerminalEcho: terminal_echo USE ENTITY WORK.terminal_echo(behavTerminalEcho);

--End component instantiation
-------------------------------------------------------------------
	
BEGIN

    combi_terminalEcho: PROCESS(cur_state, rxNow, txDone)
    BEGIN
        txNow <= '0';
        rxDone <= '0';
        receivedDataFlag <= '0';
        sentDataFlag <= '0';
	     
        IF cur_state = RECEIVE_DATA AND rxNow = '1' THEN
	       dataBuffer <= rxData;
	       rxDone <= '1';
	       txData <= dataBuffer;
	       receivedDataFlag <= '1';
	    END IF;
	   IF cur_state = ECHO_DATA AND txDone = '1' THEN
	       txNow <= '1';
	       sentDataFlag <= '1';
	   END IF;
    END PROCESS;

    combi_out: PROCESS (cur_state)
    BEGIN
--       txNow <= '0';    
    
--	     IF cur_state = SEND_TX_L OR cur_state = SEND_TX_P OR --etc. THEN
--	         txNow <= '1';
--	     ELSIF cur_state = THEN
--	     END IF;
    END PROCESS;
    
    combi_byteToBCD: PROCESS (cur_state, counterA3)
    BEGIN
        IF cur_state = BYTE_TO_BCD AND counterA3 < 3 THEN
            numWordsBuffer(counterA3*4 to counterA3*4 + 3) <= dataBuffer(3 to 7);
            numWords_bcd(counterA3) <= numWordsBuffer(counterA3*4 to counterA3*4 + 3);
            counterA3 <= counterA3 + 1;
        END IF;
    END PROCESS;

    seq_state: PROCESS (clk, reset)
    BEGIN
        IF reset = '1' THEN
            cur_state <= INIT;
        ELSIF rising_edge(clk) THEN
            cur_state <= next_state;
	   END IF;
   
    END PROCESS;
  
------------------------------------------------------------------
    combi_nextState: PROCESS(cur_state, receivedDataFLag, sentDataFlag, rxData, txDone, counter3, counter7) --[other states necessary]--
    BEGIN
        CASE cur_state IS
	       WHEN INIT =>
	           next_state <= RECEIVE_DATA;
	
	       WHEN RECEIVE_DATA =>
	           IF receivedDataFlag = '1' THEN
	               next_state <= ECHO_DATA;
	           ELSE
	               next_state <= RECEIVE_DATA;
	           END IF;
	  
	       WHEN ECHO_DATA =>
	           IF sentDataFlag = '1' THEN
	               next_state <= CHECK_COMMANDS;
	           ELSE
	               next_state <= ECHO_DATA;
	           END IF;

	       WHEN CHECK_COMMANDS =>
	           IF dataBuffer = "01001100" OR dataBuffer = "01101100" THEN -- L
	               next_state <= BYTE_TO_ASCII_L;
	               counter7 <= 0;
	           ELSIF dataBuffer = "01000001" OR dataBuffer = "01100001" THEN -- A
	               next_state <= RESET_COUNT;
	           ELSIF dataBuffer = "01010000" OR dataBuffer = "01110000" THEN -- P
	               next_state <= BYTE_AND_BCD_TO_ASCII;
	           ELSE
	               next_state <= RECEIVE_DATA;
	           END IF;
	
	       WHEN BYTE_TO_ASCII_L =>
	           next_state <= RESET_COUNTER_3;
	
	       WHEN RESET_COUNTER_3 =>
	           counter7 <= counter7 + 1;
	           counter3 <= 0;
	           next_state <= SET_TX_L;
	
	       WHEN SET_TX_L =>
	           counter3 <= counter3 + 1;
	           IF txDone = '1' THEN
	               next_state <= SEND_TX_L;
	           ELSE
	               next_state <= SET_TX_L;
	           END IF;
	
	       WHEN SEND_TX_L =>
	           IF counter3 < 3 THEN
	               next_state <= SET_TX_L;
	           ELSIF counter7 < 7 THEN
	               next_state <= BYTE_TO_ASCII_L;
	           ELSE
	               next_state <= RECEIVE_DATA;
	           END IF;
	  
	
	       WHEN DONE =>
	           next_state <= INIT;
	       WHEN OTHERS =>
	           next_state <= INIT;
        END CASE;
    END PROCESS;
    
--    behavTerminalEcho: terminal_echo PORT MAP(clk,reset,rxNow,txDone,rxData,txData,txNow,rxDone);
END behavioural;